magic
tech gf180mcuD
magscale 1 5
timestamp 1702084210
<< obsm1 >>
rect 672 1538 279328 174078
<< metal2 >>
rect 69888 0 69944 400
rect 209888 0 209944 400
<< obsm2 >>
rect 854 430 279146 174067
rect 854 400 69858 430
rect 69974 400 209858 430
rect 209974 400 279146 430
<< metal3 >>
rect 279600 171696 280000 171752
rect 0 167104 400 167160
rect 279600 164416 280000 164472
rect 279600 157136 280000 157192
rect 279600 149856 280000 149912
rect 0 149520 400 149576
rect 279600 142576 280000 142632
rect 279600 135296 280000 135352
rect 0 131936 400 131992
rect 279600 128016 280000 128072
rect 279600 120736 280000 120792
rect 0 114352 400 114408
rect 279600 113456 280000 113512
rect 279600 106176 280000 106232
rect 279600 98896 280000 98952
rect 0 96768 400 96824
rect 279600 91616 280000 91672
rect 279600 84336 280000 84392
rect 0 79184 400 79240
rect 279600 77056 280000 77112
rect 279600 69776 280000 69832
rect 279600 62496 280000 62552
rect 0 61600 400 61656
rect 279600 55216 280000 55272
rect 279600 47936 280000 47992
rect 0 44016 400 44072
rect 279600 40656 280000 40712
rect 279600 33376 280000 33432
rect 0 26432 400 26488
rect 279600 26096 280000 26152
rect 279600 18816 280000 18872
rect 279600 11536 280000 11592
rect 0 8848 400 8904
rect 279600 4256 280000 4312
<< obsm3 >>
rect 400 171782 279600 174062
rect 400 171666 279570 171782
rect 400 167190 279600 171666
rect 430 167074 279600 167190
rect 400 164502 279600 167074
rect 400 164386 279570 164502
rect 400 157222 279600 164386
rect 400 157106 279570 157222
rect 400 149942 279600 157106
rect 400 149826 279570 149942
rect 400 149606 279600 149826
rect 430 149490 279600 149606
rect 400 142662 279600 149490
rect 400 142546 279570 142662
rect 400 135382 279600 142546
rect 400 135266 279570 135382
rect 400 132022 279600 135266
rect 430 131906 279600 132022
rect 400 128102 279600 131906
rect 400 127986 279570 128102
rect 400 120822 279600 127986
rect 400 120706 279570 120822
rect 400 114438 279600 120706
rect 430 114322 279600 114438
rect 400 113542 279600 114322
rect 400 113426 279570 113542
rect 400 106262 279600 113426
rect 400 106146 279570 106262
rect 400 98982 279600 106146
rect 400 98866 279570 98982
rect 400 96854 279600 98866
rect 430 96738 279600 96854
rect 400 91702 279600 96738
rect 400 91586 279570 91702
rect 400 84422 279600 91586
rect 400 84306 279570 84422
rect 400 79270 279600 84306
rect 430 79154 279600 79270
rect 400 77142 279600 79154
rect 400 77026 279570 77142
rect 400 69862 279600 77026
rect 400 69746 279570 69862
rect 400 62582 279600 69746
rect 400 62466 279570 62582
rect 400 61686 279600 62466
rect 430 61570 279600 61686
rect 400 55302 279600 61570
rect 400 55186 279570 55302
rect 400 48022 279600 55186
rect 400 47906 279570 48022
rect 400 44102 279600 47906
rect 430 43986 279600 44102
rect 400 40742 279600 43986
rect 400 40626 279570 40742
rect 400 33462 279600 40626
rect 400 33346 279570 33462
rect 400 26518 279600 33346
rect 430 26402 279600 26518
rect 400 26182 279600 26402
rect 400 26066 279570 26182
rect 400 18902 279600 26066
rect 400 18786 279570 18902
rect 400 11622 279600 18786
rect 400 11506 279570 11622
rect 400 8934 279600 11506
rect 430 8818 279600 8934
rect 400 4342 279600 8818
rect 400 4226 279570 4342
rect 400 1554 279600 4226
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< labels >>
rlabel metal3 s 279600 4256 280000 4312 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 96768 400 96824 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 79184 400 79240 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 61600 400 61656 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 44016 400 44072 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 26432 400 26488 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 8848 400 8904 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 279600 26096 280000 26152 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 279600 47936 280000 47992 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 279600 69776 280000 69832 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 279600 91616 280000 91672 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 279600 113456 280000 113512 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 279600 135296 280000 135352 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 279600 157136 280000 157192 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 167104 400 167160 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 114352 400 114408 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 279600 18816 280000 18872 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 279600 40656 280000 40712 6 io_oeb[1]
port 18 nsew signal output
rlabel metal3 s 279600 62496 280000 62552 6 io_oeb[2]
port 19 nsew signal output
rlabel metal3 s 279600 84336 280000 84392 6 io_oeb[3]
port 20 nsew signal output
rlabel metal3 s 279600 106176 280000 106232 6 io_oeb[4]
port 21 nsew signal output
rlabel metal3 s 279600 128016 280000 128072 6 io_oeb[5]
port 22 nsew signal output
rlabel metal3 s 279600 149856 280000 149912 6 io_oeb[6]
port 23 nsew signal output
rlabel metal3 s 279600 171696 280000 171752 6 io_oeb[7]
port 24 nsew signal output
rlabel metal3 s 0 131936 400 131992 6 io_oeb[8]
port 25 nsew signal output
rlabel metal3 s 279600 11536 280000 11592 6 io_out[0]
port 26 nsew signal output
rlabel metal3 s 279600 33376 280000 33432 6 io_out[1]
port 27 nsew signal output
rlabel metal3 s 279600 55216 280000 55272 6 io_out[2]
port 28 nsew signal output
rlabel metal3 s 279600 77056 280000 77112 6 io_out[3]
port 29 nsew signal output
rlabel metal3 s 279600 98896 280000 98952 6 io_out[4]
port 30 nsew signal output
rlabel metal3 s 279600 120736 280000 120792 6 io_out[5]
port 31 nsew signal output
rlabel metal3 s 279600 142576 280000 142632 6 io_out[6]
port 32 nsew signal output
rlabel metal3 s 279600 164416 280000 164472 6 io_out[7]
port 33 nsew signal output
rlabel metal3 s 0 149520 400 149576 6 io_out[8]
port 34 nsew signal output
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 35 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 36 nsew ground bidirectional
rlabel metal2 s 69888 0 69944 400 6 wb_clk_i
port 37 nsew signal input
rlabel metal2 s 209888 0 209944 400 6 wb_rst_i
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15418618
string GDS_FILE /home/antonio/Desktop/caravel_user_project/openlane/user_proj_example/runs/23_12_09_01_06/results/signoff/user_proj_example.magic.gds
string GDS_START 245392
<< end >>

